// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
Hsch4/Mi4ypgr9UfcsEnqJI++Tr332DuuEfmJRyjZZXjwj5G8Pfray1PCi/ogbCFSKDk1iaRqZgL
s2vDFLa/YOv7Z75cgnsEJ1smH8m2KCNkP57BmNXhoKzv00zI79ZSczOvPKmNe2s2yDCl+NYbtVhD
foj5Qj0x96B2pR/pE3SOXUT3uhyDE37aUmZgiHICW6WHY06wjnJ3Q4LTiNOj+qSz1QDx9y/k23UZ
XmelNRbJVNIHdIC3SG9VVvGOB4cRwL2T3DP4acyIRNoBa0xZmXVw+Nr9MV+S7NazhwUlZAhsQn17
WvD8WvOjZ4MMr1esDdRdy/MHx1pMLqyBzIsM5Q==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 5760)
+dLW35042ot+jQZJLzFwasnDXFjNA7NeIi6+vURakpYDfc0WH3lFFp+v7tutYYlrqiACww5iu3O7
biq0gHKJneKF9xbvGP82roN2q0EuTw+H4M8u4NkSNIijhY3okF1470GneE1S4YHWMDE971Rgjmac
gbDX1Yn0BBjfVze4IO+52NeN67zB0S3vkMK9ZfNUrlGxZjt5RYH1qNsm5IMdbVbGEGo51cohh/iQ
RlgokA4e4aW1RkAKkJ2OdCTVSoGbGRBFZn52xvnpvC4Qh31q7d/FMDbTleSbp7IrsEStRdWCZwhA
FhL1RvarjxU3cW2xaQIFt6GPpUbZc0rWH1inLA3mlc1rHGJrX3Yreu8njrzFSk/4Dc6WHIhoTejE
fAtpJ/JCOhoKkEFvIxqJ5cgCZlnVofSpl+sq3VuCZxOWZ9RgPSNw66do3L11PLWLdWDNM250dyoD
MiZP4sKufJUHxuaTeKvjvlA36vsDblhih067SZaFxxkYOJeesEjlnrbhFims1OMAr3ibp7QewQwY
vSYpaEFHNticCtT+v+7au0E5kzuK7UjwzZd1CDnSR55LeYoFwTYaLciOeohe3UlmwlIMosMI+oQ1
Pv7znpLX7TtbjkexmmKl4dzQTxXOQIAeWioQdtlh9dvsnZyc/L3Rsqj+sWEDoXIxogL2zuhmeO9U
chYoosdvkuWTYhGVtHm1wLPLPnBOsAT/EXRb4aLDyBbjLWPDluCifhlIgiWX5uf6JNvfkuJZvpca
ifQnY7DbTXPVLqagU7nLRfXaWCuQDujd+qqErtnF1fpYpiN1b7H3xg9RueeFO7EaZcveV4UJWcMT
KVCxudMowc1GEC0H0f9J5AA9NiSxf2vUlwd8RJ6cApLIUYRx5DEf15fOto+NGvouWUaLfAmEP8NP
KIDDFiPETpmi9b/sgxuoVTKUYtyZ1gykc+e1fy9J0E+TiAmmTnykVv/xqWSIZ2XVKp2LtOUpEU+i
xGGZwhJAiexrtYw8VSwf/NG0nUpHI59vxc4vVwjY3niequceaCjT+21Xb2iexz/VHMTcGADgWZ9B
fUiTTf+hhk30Dq/PGNJR26qvJwCLC5m80te1BTHbXNb16LLohPztBW8/1065JkmCFWaHcvSwOLGG
c8AEVt1+p/0KgaAR6EmCGKtBFkmO6jvDI+GqIdWvFV/H+NOWvjlIlgc7LWL/fa8rfb6MLYQpe2Vo
NVyBv5nt81PyjhKESRUcCkku0CVYr8Q2DQ0vdPFDb5uikW6IbfKwFUdcIsuH5gfkrV45qBOn5IzO
8AyNVyFcuKIYJAXWN1tTn6e/5/B5rC6a8BE5ZDeHg9lMn6u3aIsDc/td7O+KDzOltOs5Tp/QqV91
BpoTsRTi38DSIorE+CmYEk3MPbrypwQWEUk6wP3n8AeILz4EgxTLI3ZKZiPpWh2m4e/AabA5rbRR
DT5uGPAK7b083qwnNqJMcEy/mpwUqh18ydS8lT+f14HEEb7RpTeUrViacx1YKYdYdv6ymmPYmdyU
0RxUjjbRO51fT1yBCvlvnEXCf/YDIRTUb7qcTzuBroOP/RiIAW8giW3RBf/USj89j+Xent/xz6Vq
zsEgN5kH/1irFWGot9lU7/9MvGTsO2nc04c1iTqoIbTDhmQhxPeuwB33sIAyuG7LvCtuP5VsQGRB
UvX6metsjMmINZneEJkIRRkfA5xsvfmFcAyFgqMfJYOlRDLpSodYS8ERZ4orY9KRyqBhl7nav5G5
xNDpjgjzavy/TVQzPsc2Jr1dKk8mTTkrg+OSo/CMHlICQD3CGpuGCKY2pQoz5HY/zBZBTmjuMe57
zaXAD7jnnHwLFo8sMWp3fSSDLpko2XSJOuNybqWMXdRPr9H8RSGJLmimZZvPQ2gLlgR67Py2FusR
dtoxmUUxb5IomkVJmUmdIBhGaBDWrN1BJ+74oJoTIteCybMGQK5vEaLZDLwmN2MfHnbRKGO/ydcc
Pv4R4hwqIs0cDCJJqk4lItIU5tYnIclSan7hkSgzW/tLeCxikYFOiBQfcWeXDNLjV9MjFm79eydG
Rd83OcIPxj035p8Cy6V04HcU9ZIMrw3c/24tG0flF9R2RxsgQrmbuWMwGtqbYokniFGV8EglUBDA
Jvlfnn1qei3yN9wzopgjuORXwFG5vm3KuLUQ85ssdR9wW81AtuHme7P++4GRDX/8iaYjlWnDaXWZ
oxwRwHBnIBTABCmYT52leLjFn8iaglEHRKWH4GDSEYVYMKhDsTiB2T9UWW7y3JGa4Zou2prGymXA
jkTqn9vYcuAoN1rgtYEJhBLs9ZUWFfubPkyuhl+sY4Her1Ek+8a+4cncplT8BH3V72f5Ebig3s9W
NY7WwX/gHTm43vg24P92g9GV5hyXbeK5kMjYwVI7VDqZbJk05G8aoCFfQseblGvNtXZCPRdlxelk
SoE3c/SZCjz6ofbr6zpjRckrT3wAwGbJ6RwY4/Zu6m0xWOVdVljvXsfvGYxd7icPzE4EL0p6F+jG
XBcS34vVFZXZr5fB/uh7f53XbKchxbBkungnrFwmnwpOKoDkgtPZ5KZbYLOh8PKrwfD2z+CclDr0
ZbsNOP915fPxG1Ntdib+/D8G7xmJW2jucWgy1XZwJhPCOZbyX2+Cqo8qmZgbOZUUq8K2ci72CSQ0
bi/rNccyAyOHKphtg73mDq+UnoWRWVNKeuqzjxAwC4ClTdeLhPgXobdiyVblzAVx+KSLKK8D795e
mVnKdB9AUcq02xbroSuJnz14DDOevtJxbhfkF1EcS4tDYn3rkgyvYA2WKGIReofEr+MrgIrpxIii
IdfaO7W7dkB2DdXlj+GeItLNMduNJDKZFofm8kpWKqQXNvrxJRWgLATI94dM7nkYpaQ84fC1hrHu
UltmVwoRiKSn85CDlLV7p5ViyxR13e+OF1xtQ7k6hBnCYJhxp//DmB3J9u6ytltY6hBraRCHZlUl
AwDB9P3Wa95Y4fsOD49heVANitk4hzAhFMlZPM3RCFuRSDSUppDrACcGrvHZ/niqh28LJRz/r1+s
zdak53MxmxTs0y+3S3IdohyVIn03hixF+yNBvkVbOVw/GmvGiSoedU+QrJattsy5JtssZ5vIcNmf
r5EpqXtHMAFighBOeWCNNkbWkOxXyMrMLR5WgZhHaA4PkaIfU00H53sFssOdZTOeeXpu7vXcs7hP
nGHp/Os4KA11Ugw/+DyuCorAquKWJVPh15OJikB3W2c5vRMocIDXDY5IsXsm1AlnBZ2wHG+eId1i
HyibMVA5y1SCUUmTM5jEkZpx6+y/3wZfdNCKuQothP2ziNtxG7J97HZSIQGnayGpJAgfFo6zo+sw
ZuwqP4BHsYx2JPb10SWXk09nP06+PJw7QrAW5QXhoUasGfYZL4nQIyoQkvHcxEKdjg0jbToS4sJh
A83awNN3KxmgBUvMnuGqWcGVjYcvE2emldFnW5UfHhTpfIAkM59lcVpwfxcAGRBlgx4Kistb4fRH
173Ytu+0TpHTh3YMs3BYksiOMKt82YQ0cXOSj2gkBPejpTPPPiy8YBwGlez95mssXsVram8+59oV
UKxnmDN4rse9IyzhGsdovTMsXlkPKG2Gc0sTE1MNrLVkXq8jg59eZVr7sb+X8JVZn6aSTO34UMCW
Y5zjJpMZnRfcUUhfjEBl0p4ABUcybkPEWvGzAFAZN7fTMJWlF1vBKETSGfpj4P7HZlwsIgt4Vw9c
irfc5Y637Ai53BMqDk8gbzioUpxYwqqxu6Fmuhw1mivajTCilEE+D9zq4ChlFKfn8fMp9yIxjqow
P8P7hO2D0LMTzwNQcTPMazicLqOFh/WQ43vWJi+5YQFJgTwjKvneOIsw9TdKRN/XdnvqWJ2yc/QC
6s2u5aMQIR7zJzUDudWEYoRTQOVPvW9jVOTNBCn28JxQwUt6cI9L/EJrL83QLMzJxA+/cXjBCifj
AUiP8//Ii8A7NEjWAID1G2iphrixRlJM2Ad61ppo3c2TfpQzlK78M0CSHJtYQBfSUYxypO5ekPe5
kiAqxGt7sk0Xe3fvZ4weXSTCehvoji7XliGegBhv97Yr6QXV2HjubEB+Ga059Ua+cihypvbx2uHw
+t2VxrtfsY1bC0ls1lB7Jei4VsuF+YulYcDE197tKVuf+c2vYO/OzIaNQ9boxhW+GGhHB9Qz24tv
8VwUIX5RhQkzelVr4WTZFC6gYzEQviKGKYqh6rVMd3/17UgZZhGzFvA2+MO5ZNSoEbSPA8x1hCJD
W66lezemAnPdx30jZssIU5clpPtwIPbBH1cNcqu1F9jfdb7e8Zko+z9s+V431cmkROx/hMN8QrRa
aujc0LUQYItcFAuVgjcDltncG70p2ReiD+SJvySdkFII1fmWZTfeEtnGGUwzMbMSJxu0e5s/tx0M
gscdlmux2/w/kQZUQLH8unDpciVV5HYINQVfNmfdA1HIaTnxBeIz2JBzUfB+xoY/nisvDOtLGSzW
05ipau19ju2QVrXaHI7d4i+6r6jI3f4uO9baVSdDkK0lSD+jux+lDqanfllfs5BbB4jIYpUPsjlq
3KRdUWP5vjvTZrZzQCtTC13MBS4O/F2tfVac5UkLJJ//bOc1UHp0xbvEN19kIP2eer89e3dt3mkm
jVXaRecwLINy4JQJRPkroh3zReViyzpzwX9IAVR7cuQT448RXe0nM7j5lyoPBxjsegE2QL0ZDXIz
S/gjqG9o5o1tBR324QTTps5ClZnkvkn9UmG3HOk7dAYSQEpWlkGh7YMvMj7qVPUIj277GF77ryHS
lcrawbgn+JP4n4p3EGLJ6ly1tXZtKIPQXKGkAGVjsQzzAFus7OIATle8rAyTHPrB+DG1p7bbtUYq
fwLfTJLhVniRcjTgxtPplaFqXly15umaR7l716O0KrbNNEZsMC87eJWvP13ZhJOfXwgJC32e4NyF
8FOR4T7x3aooWbivsDbEzDXZMCAUWyx23qAuhZhQNBDWOBskjcdlVB5Im5+tzKpyWGdOobzQrIp1
RKkd/dGhKBzFrhXRz+LT7BRc2enpgKUFWyKr3t0ZW39wAWd+PxFOYI5Ty0NhhYH3SFTnpPcqILUT
VNR7sHpfgV8+d0VsQ7HcU1dLpa7X/emJDyy2rUhZyq3cMHEUm6kgARZQcdKV2GjlbYevwYe/MWiD
T49E0sAo3hDnBTbX5w494duXHOOKwOh8FW+PWfKTBMxNar69WLIGTE7ZPXqDwukumM+OIuo/Is+r
j1sOhTu7OgQp4XNQ85WtGaz3L9KBLTJ0ALx0IzRzFsIch3UZbZFkp2d5IyiaT2UGc3M2FwRLhs3S
osBsQ7jbPOxE9JmOJTdCPGdoP9gKDBjQs5O2DGBxK1ZYuHZcR6K+nevKzPna3Tl+LDk/Dsq1Le8n
jeWHmND/ec8x5xRmvTglkE+HnrZnbIp4i3QMEVVubawjWvoDzZs7KJDsnjv8GOJAxU2SjeoQ3SE/
xoO+1h06cSAtjEHtoZiSitIvmDjERVun9+AlJ7zP/fEC598S7Pra7CUxuaKfSQmbJrja9+WkHaC0
ZUMe67LWpAlDZVA122iav/K74r8bd5D8IEY6lE/rqi4QBXS5csalbO7Ie6CwTMb/Lyut/zcpOuH7
UwPvfkgUvC4iay6yYQirqDNtlnUPI/lJ6ZcKngrMtaQ4DF8gQnWZDHrcbWVcTI7DzvrFrGD+TbiU
PtYmKLjDCUHrUrHBgH7ddoTRybG7e7MgFQCsSGhexDZB4pkOC/+/FbH/tEVzYTZZR5lP0AN0NZta
VulfmexuiqAbxHP+njdR14o/24JNAom2yLWqpFo8fCSXoNGgEDx17uNvfi3/wm4kDmYK2xZMSbTC
SJhRlzL8qbwN5vwuJalkwGfnTFkOKwcXzgjPmFrEMHFEjK5Ag4BDi5O+taFIjUzZe/V9XrWN+mKE
BV9qNa5BnSie0TEFlc4+6TK8dYPrjKdhVBE5EvAfXPtfQzkPLbeiAzxp8Avlro6v/TV1slh0ZaeN
7hq+auzwV+Jj3Ss9m/ux/DVZm5RQ5k3EDM6dRObokVns/OJ1nndPeIc4J9GiA3RuzlKiphFHVFh+
XlJOJ/2Nt2Wdbtv6EQHkl6wQs0zUz6u/bCGYSzgpI1r248Uzb5MXxlMzyIXlpvpB+slIMADrf1Ky
QJH1/kEhqKJdmfPXhL009L5kUNyL1tNB3eo5b6zMYfKfBPiq4sSdmHmZ0ccWTLjfH/0lhexCVInp
XG+enGvLUlVFkBY9kU6+wO6UpDWLA5U2XFWcJ05jjBFE74YJb+1gBpv30sQTEnPQjs6gJjpkZ8fu
0Vls76kYc4rI121n77HMniETOA5DwoBVlGCMIOwACP5o5JzZgmevpNn65PfuXYKpa2wknI5UJTYN
msJifnAOT26u4tSiP0OFrKrzxvPV0ZMygsy98empRC+T/rRndzGDSrSAvKpOjFOco68iYkiIidEr
rO6es85Xq/hqpMXF7KPnlOMMH3G6nBCtSsSOOOrSvl1Kqhb7/KT3YaUTZH7VwtFtDm6D6hib5pp8
gA9fjqV1aLReBB2LFvnp70sFaO1OKs9ksaAESrLfzGA2dLdRL26Jz1loEgx19ffGCePCunluTYhX
KCw7RU+W4UhuYq93pQVJsN6XSfnoytdQWOJKQ+edmeOCHnzpeqZSdRodU2XqM+xwn+U+2RvsNJ52
wicanU+Hz6FcSDD2tWN1iXp1EmQk+hzWtqnEy03HyngKcBD/p1vXoCEFdPOGVOKaE7cjgSB7+/PE
hBIt2KPJWyXmzAbYkMozpfL2eWoFBHKaPVF/mi6r7ZY1T4UTzqNFxGWMREcpUV1+k5/HxCQt5F38
S3A9kVgiAdWOzOnbz1xz0IM3OCbMZ3GH+jQy7QGT6TtnYJtLnEU4jhYpa3NbpIk2YZv4204noQ2T
HViZWsUvbOmGpYI4ofKIZC2dt8rT1iz77q1VzC08das4dLSP0moxb6FyrZou9XSCMYO7E0bj8785
ucOOAEeJHb3GhZqrr5AaJQXd20HTUI3xRBxeQoj8aHpH64i42Aufv6f1JwrD5jvHTcqEje/1Mjuc
Wz26vCSjHWe9TouqMQR6fMNE+aZkaIq+ProxAvGEW7cOxQSLDth08mGBSyYH8t9Coix3fXiNLf5e
YL42PfnauRgYumndOErlgsh0S5BPeuhMkNbX7iYoNRRJV3jWLsXZkhEzjgD89r0ygyEfDfe//HVd
C8UTYLHKK3o2r21ldoJwt9ENZGM7qFIJGGp0byEPC0GvO7WGvvlFpwaxKcMCdPBOJkUnBm362sUy
WXU+EKV5v7TC99ZLUedHtuxtSA6cn90+D6H3nSQ9Kh+ovQfI60OEMQccnwOPlNfUqa7ZCV8V+/fX
+2MNMYH0kQiwccHcvqV47E4v3XzcqKQepa4RX+tp0cVr1IXRMoCFVEHt/NuuUrVJb2xs9ovvS9PH
QwXcxVMD/UIL8/esQrgTcwxIwYQGpyMXGb8dhxPCxESnv6VlZ1HmWMERXZpek8gasZYvHpPAs5AW
t3FiQI8Em+CXJnCoKdVYfjcS4XCnoUPHfBJRcoqeLQpMZ2aBpcF8U5yPb8gN1w9MRfaknaKl9wHr
72y/G+VrJ2ME67gWsATHWRSFD/rgarltGwG6VUloP20hNG2R61kIs383TKaCUAl2U6Qh32WnkDs8
ZD0N
`pragma protect end_protected
