// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:38:09 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
UQtxXTh6stZoP07ymn9R0q0nzJdCKI3jGnZlo1ab3Yajq7vYOoHz9mulyHMPiPII
ct4t9uWvrGAYtPEgBOYWjNjPvEQTZ4aliQi2QF/MwvOyiq0WbeKI61j8pST47rTq
VAmMbwuSVZmeDIGjSv3Rf1zDWtnkkBIV+ETQEyydW3Q=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5840)
klZhMwGluAFOsM9Y0I4GMcVqu/hwo0WzTYPMhXbdNS3n3/xF1yp6/Pd4NSznO4Wi
4XxzKwBbmp/n4Pw/NR0ZAT2bIo6kasFZq3eRaKU9Ff+7djBT2ID3p1akvQ3/3aBt
G4RkZIYoIzPZNewoH9qH08CGPL5A0dqAREH4SOivYRoxHDRXnYft79AseLeUeuKW
HDsZN+QySaC9wLKlF30odafDQsrvvwydzqEE5VGrCvYnPlHGNl4ZCIY0TR5bJpI1
peOS3jrFqUuXZLfq7g6eQh9ocaR14pf0per9+L/3q66YuCFL0OavDvkseiqoxjgY
jCF+cG1iH8G9z6bbzWx84rrCDQcQaw4ZaNh+svb8a73r4EGxOrI00FARZN10m1Tu
V5rcPcpi3qPefsVft3mEt9zQ0Bus8ueROls8aLh+aNySe6ppIu8aQbsI1BPdkIvf
0gkbbMydRUIcNMiN5FmM4LZHzZfVMT0bh6Vah4ugi66DGVMkHYqjprKxFVBZ9Hzn
KXgmfxZIE2Uw2esBZedxcipCGXTZ8lwY/EDP3fBp0L7spg15aK6k1gsyk2GI8w0K
yiOSAsUG/cX5QmKCV0ZqcJKhKRdduYNtV6UH9wh+GePJGgwmvhIPSREcQ962YsUE
AXHD05nGRrGU9YztDP/ILWXLbokWp9Q2hKSEKeU78o2bV+Sdnb0UXu0mrJx5by8k
FHqJNSxWY9Udw7LLrUpnxRkMCePl7nT9cDNXmhbnD7QH5Y+jcbEJKWrMN2sdvnRk
HtUJ3VRPLzlCi2+Uyc53Sq+8aaAQpPcAl5f6Vu9HvRRcFFN7zSEpvtsx2gFIOuHv
YmVwppZYkoECYlfJd7iDIg/QpqXp4HbQBJ813TxvOf6Ho6zKIwb3u/fchd2jlBXk
2KVr5tdHMRcwxATTWXpKtvLfwG+ZzFXnQSnUm23kY2EqtY9Bk/sm3bNLtniSdWqb
1Yv0QVDpPET6CwIc94C1+rsSHIQT1S1RlNtdC/HQ4WrXLtr2TMetJzBPq3Z9EuyU
xWQ8XT9eGn9wFdqZFscrjwsiwKqa8BtqkdZ/wXFKfnrgJG/yswBbRYWVJmOjwsEL
h+uKGQS4SbFhjxV13gRkdav1xmhnc0UOCDwxpoJw6FB5x5THQNOVC8gA0qj56bdx
z2Tr9tHpt+ScAwr6GmxOG0pH6gRt0jKyOxob27fodcPxQBtIffPI95NMpFYp5DAz
CU9m273OSnUC09609Oj61uv1I87Fv7if5JndZdy1yhV0ODhlxDjbq4W0xFmEWm0F
zmu2ySlsLFiR1K+3Y7R5QmtGBsYt99Z9HitnLHQ+z7CiI12cZZd5zc5YJw3YVYxA
7TlYMTvVbEVAK7MBFS0+pppanJUwLLxqt2YOIbCvRt4S8Lvc54MTtgFsKkpq2NDs
k82+5X9fP78ag3TbRHrQO4k6j4dbWl7iMPItZ15j4SFiUjameaviRObTE4IkK164
EVEGAxgZDhiFg6Sx9/FdBDAO2aUxmNEuDStuse5IhxWXncfFsjw/Yx/Z8bcWHYGx
bP5hyW5Mh3BM7RdN59HrwOVAefDiQ841s8yPzcKaQz4qkJ1YsufFHpPJ4ZSc8ZR5
GyKZQh41jIWF8ikdbpmXsI3DAZ0S1qGIVI/Hf7LktT0+ESLzMftffdB4HMTl5hnT
LKhGetmGl2u3UdjIe91bXY8oIaFv4enOLp4ry0WPvRDvhIJrq1uq6LczAuSJUPBh
248dRP4SdvoXj1yzsliwFdE1/AtklHy+7ByXxDkSuZULGF9bz09vfXdZpoiJrlQq
mRFGq1D37YAn2W0Br62Smoe5VihTq9zS71oGdSoGDkrZMlc2wpLFGxjEfUZ6nOuX
PtFjOAhfD9Qa6az8N8S8/AUQdGZeay3cTbCv832Toqm6kY2obTeIoexShTcAyeDp
Hlpgec/m9IRLzL5EDAkdrSkJdN9uxY/Hl2wIDQiX38GRTP9vQdy7ZpNxiJNNqmIY
K+XwK09CwuK/jDsAAfI6aK8yYAKJVbnHxJQ2BCUQtX9gNDfL4AVxCsf6ML8TmqA9
R5Viu1ofL0uKolJLrnoi6NONpHp2Vt0Tt8Nmsq4Inx405xEiAl7zid5rdoylnzWb
mKHHbl/A1/BzqUcq7UzVOFQl+dxGLzs9x4tQ6ZLjhoEmsAYhBO72XBLOKVxK+pGT
/6Os+oPUesOXr1Vziq1dvufhoGPh1O4Yds3W0qs1ZNlZzbWov2FBFN9wuAwgVCNr
LVWIfdHlWw/oMPWG1GuVYET0/s6MjQM1u0U+wFx1TtGpixuzCd5H98tVIBcYkkaZ
li6QL4yo5GO5zAoo7QpymP6i+rYP5CSyz+N/tgguhEHTLYC3Qe2gkDYn8k49xElB
cG3OYrKeeQdvYcRkPdlDXN0G5uu3GVg8lfRNrSuKxOpYMg3UlfeHu8Tt7d2OfsGP
0Vym98rDhQaS/+hCGf48QYROX4h/WflSceZEwzq5uheXNYwrAa7nCAwYHfiIUQ7F
P8mSP0LtQvx7VEQaZLLq/5rFz/M0Qc0r0eIzV/5+xtlxF/xRW7MthaGtmix4F8ub
4GtcmGKFpqDtCFpm1cI2igigy+pw+v7zQ3t8mYhaNj1PNRYsz1WnCQsraQ3yvW+M
aIW55LBdO1z6oL4JoJ0InvrykzK7mkZItdCZprvH6Y+N1yqr//owUPKXXcqE/BP/
T3R1S674MOuKOmmBfwWdmdM/kdnlmAql0re5hWkODC2y1sza0seisOdgkO57WxFN
Q0Wd+1vjAQAJ27R7P1upPzSirbp9sQDuvYug/2U5MvnnNnuF8dn5hlDhvzzur5yB
/Vt3xASVS1/xBg53SR0Ckq1T0ofLcWOrjhZgED4seDtDAUroYbTUNe0RQS2Cy9rL
5eVYGFruEX5XILvPb4pJIbpAot4UZWqCFKFJFiC/7uV7dGRLFGNc0vu2q4Ai5r49
d6dGW0OZytsN3ZCmnVdc8hAaESI7lsY99UUMQd8p7NDfnY/YPgmcqOGsg3EAKctv
8GspCVTKtKIuBJXwv3tfgVuq3OoXlNSlYW0gY2LpruoJVqZUx/irgM1TDNPCyHK6
pB0lDuciMRcCuqHnRhiTv5PQzMVH/THBj8gTF5buvSdQ1nKjgocXX7BSuM9/E3MW
eoZUpflQ9vk3tmEqtmAL36Bb2jbll4dsH1AP83iyUlxWTo+gamXftp5chlqJrq4b
Yzkq3H/x8BWtiPZ8nKZsg7OqtKl9j/Xp/hlK/1Lgh8K/E3zOfgCFgyE97MY6d8xY
eZm8JjzJ+ieOc3qrktenKTX/rhx+owfpRebbPhJ1cMtCWMaKo+XqpuLWkEpHLX9m
yb+xl1tX1+a420k6Vf5sy0PqXndKM5gFZ2XU8BnAfJjJbkIfEru51lRfHmbaewNU
hVuBCQKKbLJ053eVsAovzVG8RvW/SIHvt2SsL9qOIqH1LzF0K477R3fh5RCM2zu3
bTSIOIeXUIgOUtA89ruJKHbYtROQBjHaMlfZJarIDYItpt+btAc8y3/EItKvdXKE
gRQA0fkX6OP0WmVc6+5hV42pZvT9gTQXPiCDV1nG+TqqJTkz7RiDcBbZcZEpFXQ2
FQlXvmRiG7fEkqHzYv9MEjwAwtYL/2tpYyWeDHEsns6NO0p6q6h0S3/l/xmsGfJA
cLeugLesRfLIv2z2kU4oOwZJ/QAkhGlYU0PRZNRnNBksUv5mm3rNp8u2DaXzr9EU
3QqhvrYhT6qmCAmULeRIfZ2+TShiqG32u5dKnb30eiAQCqG/UU9vHVaN9yQZJ1fT
gSDyiyni5SjOIOF8HBj0gb6bpmrfOeBzWjHY9rQahIIXjBMDLuA4Tt+mU++umT47
WBSKANGnPQjWwcaPbxsoMvGmlbKQAh12LCVanVBeYuzJHiJg6zaWIWjiUrwqL1DG
HkxcU1zEuTU/GMItXlPZ8wMlRJxvfGoFkq7jbf9392+71J5Z/aEpUzPBimZv/fSj
Hdq4MAqTSGvWeFBD2/zaK0pd7UObYXpb9gl30pvnBxGJ83oo+KERKMoHUlJpF/qg
tk2gj3gvX6dPSLKhJwFaky+feFJaDjvHpQCY0M4FOxDTLcJXtcfKuI3hcoCrWerD
0O2dDmdj4FcOlu9N7REnnHu7zk4aK73nh+9ZR0HzskLA4zXEbGij+QcpIX6VwCuq
xMnRgTy825DWjt/h6q/B5b7QHHdwZtzTShXnqGMJhSTrlC52AfXd1XbYVh7YXKaa
DVFehbYzzQyKFPQnwKxRz8w1UNIqT7P13Ny57C1Y/D8Mqnh/LkoX6cgqPe2oWZWc
DQMIdDtQNlTk+vNpdl9Kee01v1iTUmC1ya++YdsUXIApfvi+lLHJPRYLkIhuNnW8
/80Nxiy1g8n9XA//mFPDM88Ao/b2sD+A3wWWUNmmVnCAxs7NrQRqeRL6pshxPAce
I6bchCdgwB1sIX0dLq7HhaugFjKisHPLY1U//JX3Bw4IWGtTH0jEXRGaA+wB5eKc
fWnuLKMw4z1ZOnVnEYiZJNlbLC0aHs5SKYpvM+L2Epkrjg4tuhnTH2hNnd81XLrt
WqxpG8UPdJ0YeauqtdERlw80kMqG5E6I/Oj9Yf2j/DyWp5N1JAc3PJIpQS0zt3R7
CC4ZwAHchknBC0Mhglm7Hcco5WfaSQLzU2W1kjkqyH8Fpt0fW5fXvvJMgtLVv8Mm
IpaUFMMRIu4ygz3TleDKOATGJAaNyQuqnmTFd0E2uV5q/bvQZoU9t9aDIAelf81+
39lE8oTAMeR7kBEA8oJeHcQS6OQNbMqJbOyomPSi3Yf0ldSAEamHaOEkstVpmYOh
I7MxdwnqWdOpzSIohDZdiR/vqW3poFhx6W3P1GTd4zC0mVlNLj9KBwwazWguzMvx
edQ7+c65bKmMyxgEp4KFPfIv/EjSaxLFyvLX8jW1HceYgcU9idJ+59ZoB8j1TjU1
VkS+TcnUXtTMcK/MHXagAgdpxAPNDmrRxM2T8oW8OpGsxkHPbVjxc3lJXYjbfihO
gsTXeP113F1BtSzH5cEWS36Y5EPArtBNP0Av5YbQYTNNoE0D8jLLGEBMvxLp1dPe
Sl943PNc3ekq1vAzTqXgzVC02nHxs9xJAcbwu++y7IoNG8CjO/HM5kHX2mgTe84w
3+ZftFJIdjjtW/8BbGou03aj6RPhjnjqX/DOfUykHNriHjZ1txQVwwbK1kIQunBY
Y9aDEfCdDZnjyt/wAZF4I21NJkmu2J7Ua2MYBMZfWTNUqZdJR1S4UTifuDDwJlDY
xCf6azwO7ImM6ChchQNqD/NsN9Xv5ZgMykWgK8pHZX9EFto1IWCGuSvCiG17f/S7
xVEWffol0sv2Pdc0bXCgTIv0wBzzI+K5a+Eu/CS1ZLW4DHhfczZFpE5oJTccMHmO
38bKUsSR9oV275H9dkuWB8yRsEFrDvbi148es12xr4Fc7nYITMRhg2vn+fcuB/iy
dVkO5KxJYd7zJ/vYIa/gOlA41yJgG7GYCk9ACXThKI5n+RRT4HWBuFr+ZIfwme1E
cNZX6LHwOqvAm98pkbDypk5AcpVTwh/UgDSxo6kIvicYRl1s9aZjqJ9qiIqIJhbD
s0wvMV1+oc/S9ZgRCSbMp/pPHE6lIM8tYW2V4Ksr2mq4v+i/rtwcFtbUGPBbBmyp
2x3Ox16Jr6GM/YqYtUjGhTbltuMLj53RrM/+U780Oxx6VxTJt6vGs0Y3rJnY8ud0
QEa/PfOBxReYTr7O82KaMgcQbvMA5tAGqNc2j6JRygXgdJKLlW3VJ2Jwqmvctm7O
7LJ1aba9alVpSaoS1QhCx7fqCJjqY6qvD1KHHKKTOac9kQKLCru63/CazTC/0Ahz
LSWYjOb2yyrhnrC+zvjEiRM7CH72nHFQJ68AICEH1Bkx+cwsax83uLG+M39KYif+
QVPFnRn+uzvcSWsWVVpCVJaOnJQZnrDla2JQvqWBzFdMHhOJOlZcOuqA1ibUGrnE
WSj27oHNYBz+ESePiewtjN+ZLJ1B4pszIjh9oXQ62nhtjRTwCt0dynsdsYzhrWUF
COnhMMbX2RglIwV7xI5gMkb3YteKdheUvzNnLN5PSPjkb7cudEgYC4WyUpG5CFTo
ctnkmWOjAvVncpEnvnXno/AiUouZqHOCxiuTePInZvWT2jYqqkxpMqJBc7KI6qAR
5NErvwg7I64y8cqD5wMW4/+0aAtc3a3UaqmM6yjaG+gGjDGPLcaoIbvoNSq+NR/N
dR6zNf42VQZNdwhKxeepywyfI2qPJ30Q33vLTfmYhOel0/nb3/Lt9850uGaqU1Us
5ul6yYgGmk4nAvuBVBJI73Cb0vGBTgmIyxOgOi5uJVIRU2s9GHC2lNcUR5JPn3FE
asaFcxVUZL/6L96ENNFJUA/0sEpvW8KqgYqcDriVScXogr49MQIXjselVoV2C+rc
a3Y4gknJatsSH/Xgh6tMb0JJBP7ac+8mBcSUq/ili/932Iow1hSmJ+USUiX06Lhk
6jWZrwLxabUxhgOY6ZKfD4lYB0xnOmM7OmxwHLAXxtIwdFz4Q4kjvS8eUNhL2cP3
Yd3FjW5/6HPEH5CS1uHoddlbciOCG8joC5oguQfFeuCn488ENKAJWbvex9+SE84O
N0CumF1QJnNUCVKNTkU19U7KPC2JslySmV/Nc4GU0INoH2oz2PYVWwnv1wvJb7AO
Gj633fz0euuix9abnT/ZmP+G77V+7WkenJ+Md+hFrTUWOovkezh9omHk67PkonUH
x7vQjkh7Oc8D9QsCjFEIOpZIN1WzTI8IH5hnUjgQyBKvK0bydmha11a8okdf7PhS
DvmUc3Kb9EpoJw/9ClEATKCK8R5GUa8L9jbI+aUEB0w1fe9Yr06w6rZWX6EfrEnW
8Chl9N7IQhkt5Qnp5iksVJc/fdBU8paKiTMEqfvsHr5yMLXQbOiW0Qm9iwxaJ8OB
VghZZdGkINSxb/Sv80VprbsrfOYxtHZRx1qdEngHpU02kOHBZS2LML3bFGN6Y7js
kmm2nvPlJyUVv4GsYVC1R85lvItWUv5cWp7KP9IkZdiITpLwj515LomIwByNSpKx
y/J3V5z7ZdSYiPbb85cAiT516MgEt2vePuMpJJbaIuncpysWImCKJ5F0e/NeygGB
7emcvOQIf4VYZg+2/DVsTRhCBP2jOPQGM5UMf/lKhn4JdVBeWF17GyfBd8xG0ZsF
ZcKQjlPPOnof/mDYT50haKT7gamGz7yc22QiLGZImWO7/Uwc/duCrdqxbVCFD3uN
vUVMCl09ELpTf8ElPHts7No/DQfp/59HW7ju6pWdpzwz86agxm3O085C84Sfa85r
QY/Ut0/lunHQB9zA+JjltYUYKvBDltaI0HgodrQINOzBGcWK1Frcrld+VdNGgYdT
f+jFZwx4sWtUxYXOJ5SjNyP0GYLCLxDUaWVm5vVpaRXEZK2dlu2NNxUx/cUWAtqV
RhglDDCnsM0yTWEgu1XDT/aXXGKypuDWHPsOaziX0r7cX4nxIKLUJl/RUmaoLSc+
s5oRghVauMkbAOQIowqqRjaWEbiHW18h5pH1lSwo1c+70Py7WhS5QRv9YQQAR7uI
gcA0N8ohyieZbGOT9WEdV8g4SLhNsyeV56XKU8w3lLeXBRhhLbX/ZH+g4Q3eMKtE
FJrEufWvOlx2TrnjF86f7+bwaV7Z3EFHZXT/O3IbvPGrwIUsetqwjhZ+oq+RbAF2
8zXQWOjxV02tk/2YGFJLsMTR/aKAvAEmBO83v7cPnUyf/DuQ+M9wS5l5WzgGIv1f
vzRv25t2f0+KxllkyrkBRoFgcGYzOCiw/5LaIBzVeuo=
`pragma protect end_protected
