
module fyp_clkctrl (
	inclk,
	outclk);	

	input		inclk;
	output		outclk;
endmodule
