// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 06:38:09 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
J++G4AZXJqg48cFkrHT1DBiKJSQWljymnJS6+/bSNqsA8IpbNX/o2+CCNck3v6bN
gJ0ASSvB6MJ1AQMJozeROpQDgTkGM2wrrpBAMe3C3C7n5qa286YlkpyS2lEA1Z+h
0a9+xWFAUR2CKhpD6MDhNk7/zPlE/4+GWEfq3iw6fTs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5344)
MzK9jj8hQN3OEdVJzRWu0aRvdtrUETaaWQn6ubMNzt2aMGDqojSKyeCPVskfn8TD
VOhdAhtdlJxRMgkJ0QXeBaGL8+EzznacYGecOh53Gpn/LqlSZq8C7VOsLNxsfKNH
anTeca0tBT+/BoFb/NC96UzKGB3ojSddHOeNKu1kLgxWCGEDH9zWKZhZBuuGRMo1
VNAMuqwt+Fv6FXGkQa2X0yb5E3Q55LYJfxjPfrSX5KOaDOWzruGWlJqo7627aKiK
VbS0pJWgsd10NUFeM3JhL6mZnR30tZZM9o6NDKxx5o+mjuHxfgLqNf/+oeBAIXHd
amNjrHzI2BsUXKphbDOj0EJ7dMlsaKHXWsP3hqhWy/xbPStwPRqZQeoxkMA9qT6X
k8Lm4EQJeLm0xXNkgfwDa7+o4Yw3l5bqBwP+rvrZ/oYVo4nci+mskiSjo71kXPqM
AQ39WO2SGBs39ZO43SPWMX8pX0tNINHhMtAhD1E/noUA3yvSe/eLa6SWHmJtjEnW
l42RFDzVqLNsNf/tISep44Z4nD4NEIMoEC4QXMh3iW5ELvcvkSZYbx4dG04fvEVH
UUMNJZYoE0dTBf3F0d3kHR9FmOnzoD4FG0nXFSQ3rekfOOopafUeW9GQChEbwnc7
2yt8mLpP3IlaCu8V7dsg+bXv4keRzXi4Ef26w7EEedsJIlAokapgznCV40OlP1l0
BEfP1CUzgAVNA+wQDbZEIFn6r/kDEYThKOXO7cbLEVoF81/IQhyqyE5txQc6Fnkf
LKGHwJ9DpsrCdqYuHJDcK8itJDRfu5y2u1kw59hRP0y6RXXITZPmdhe7THAm3y1k
H0nlCyxC7bcmnxbHZCfj/+pgOnG8HFOJ1FK5NXd8ggS++rsDv80J48DrvfrfR2nJ
Mvb5qGzX/TL6KogPrWPd8iJ8dQQF5kDHhnsQUCSzqk2KsvTmVTY7EcJ1z9NbPdpH
Qp+1dhpcDqwByWk8hCNZj/y7jb6PUg4FiwW76ZEsMz5s+wHrgEwf5IXtLkwpeywL
nfSSswE3kOYBFTqOtjmxccmcxOFaXPMHiKuiNnT1LLKdpFjQjO2LUu9PxOO8+y29
gc1rIhRNcobCkDekRAaJvOE/Q258vambbl5W53acPC9Xy1Nd0AQHpTCkYJzgc+nl
tfR7HQi6J5anO/ESTMtEQ2cgHquHJ78MyCBbDhtR1U9LQ8puxqSna16QgvhRT2Vy
ul3W2nfmCbTYd3fMlKrvbPkIsfv4mshRoahG5P3E0W4lwNRqNuM/uf6EIfeNRETG
DKsrHlPD0Jq/5goXqzc4LZ51QHp4l0PiOfFB0CJTxw3epcbkmYLFr0EvQ9iM2Vhk
i3x5TG5jypDjMH45ZCVafAzVbULQAc3QZ43Clv7VJJ0NPXiX3w8Bn4/fu3jGD+UG
VwTy0Vk+JgvBjm1OKnvL220dpnyYYwsoKrpyuYszKo1GOL49GBdkeX2c3K3A6VoO
xmn8fr2FTo4I7R4npTHJzsuiB4mDEHaiaFbRytAxCdD1q4wPavBpRr+LUMH3V9Qq
XkaHnK6fLzNebt9qOXtvN6ZVu+ySJMU8jLVASCnKX2f8XHfS2B67R/ryRPijYc4g
9LKJ8V82Ayh6nTYbLUtoGVWFLbO7An5gQV/puhp/A6cIaZkcHa+wryUiAXQ3/qR7
Mg+Jdtwi2p2Y39G928k8XNTvUmxTXUbQaI1IjQg7l8TMdob7e6kdy6F/FKW9YNDu
l0ves7kwnqGWRpcj2H9vKv619EpAL+nXulQKIBIel6RfamsypZWzplR6IMhEz04Q
3nG21V2fD7YJjAxCh4pAPwjVTICr25qTQ/hvzOcly4J5zHYVIOwCja8XMajAKY7r
UA9Ok3fpM9LWdo2kAUYOMV6LSZvz5oBEkdBSTv895cVv6IbAeHBPRdRrDMCLtF39
XZy2wt7u1P4w1ev4+2aWlwF6xAU76WG1LHQ0JBgb1kOC6LkCV3yPkNAAtLLwCfZS
LiyeV0z0d5YLd322dsToHjRKh4hO2q3sICMMABM1m3h2ny5SsE65wiB2zgPSGE16
1oFkvus5mQV8ghGpAMo03rAhE62juGjKy2GwSWGtG9N3IgKSJWDBVU+8opNCmU7c
NYZ8N6OlGxV2aETsDJgHRmBHMK4DXsuIAIoBYs5FRMG0PP2Yjmvpa3zkcE6wiXhM
GZ3t6VvakegL3U6ekARh5bn4XD0yEouNR1Ms7knKfR8fQhmEObZL1HsBqMQSdLmO
pI3tRy0oJwhIxb3civrP69fDVJuyyGbPGoErdxivp8ajFG4tJYeZcY71w1BDSeaH
3jmAhxhJWeZsyl9PbqalajeW6H64a4jzb7j9KDT3Yt206he6tRScda8zGT7ZzsNX
O4OGzMs2Y5X81siklUsSvOo8qJPF0caN0ZSn44oU84Lli1910w+4WyF2Pi+2e6Ph
Pn+jtFzcqUOcd1pCxiTvtyMfzKkkcHXrzAcSTQsFTxNiIXbV3nvtPl7Fq+IyeP2F
C6mF5ez7nZlIjf7VUNsnEroZUgFWACJ20cVFkXTdfaOobVhGUj1pSlu4KXoA4Idv
A1pdaRPOdI1f/Jb8PldUDwL9fEkh1SVAHcbYq6/Lr2oeIas9gx5LtiUz7aSbBvZY
Het81UlGYcZ1IW0OksRcaZbQAW/n1k3GlvqC9OyawX/ZTsH3bPvlP4hGmQ0qbGx2
IFAfC0qVoNemkw3jWoJDW6R0LlDvcL0/n3cJDLckox/k3SOdg4YKsf2zyvhXPQKn
muw1WwqmwhwluSYaJqZOdV8EoyJKbWOGP3H8e+ASFfpoexhY/R2CPWEm/e7uD3MS
yBx8YoK4wJa3p3MF21EypOv6tPfLl1XV6uYxG4bQIa69u7ak60EsxXTOfJF5x3EY
lLIRvsXWt8X/nOizHhDPwdvbF2TUBR8V9ZQ6iehcowC/+Mj6iUS9yKsGB//0dyod
mZryPjQvuPXS96PDrtij9HmPNqF6Ziz/+40uA/NB4W9prNMzqiVZlmGIqkktkqqZ
6zQAMT2OPUB1561mPaPByuki5i7hdOZ4cnN8sNAiT9RNCoIqXrGG3gUzt0c/eXv8
PF8YkV9A790ZDCvx0g3UL7ZuB5DfgwDRu/Lrq/Ui+vnBbU/RMDw++iP1EgqVmwrU
1RGPkxNYzyUK1KD0pkdsk7cSuOkQB58fPitdgW5BPXGAIobt+WK0slkka40J3lSh
Fk8sgS8hJ5Hxj8t5Yh6bkynzLQGxbBCoRzOrhZaDwHbf++y3jrDTz1EE4hzkXbzP
so3tTQWLJQDJ2ZVCUDdpRdEacYN5OnCi4mXAQ98O6COOlZ2PcSE9rvzB4X5M9G7H
TFVG1qCFN21rCG0WXIwGS9jNaBt5t4unkBD27ySi7PAAQvasTISJuBG+wjIUk8N0
A7BkJbWkOuXf9Pm4uCms7a0jWXR6aaYrehOTOMdS14D7PTbF3nhNemt82lbmF8i1
6GCWKtWUl8yyVxPMhB8tRd+/HrAdZ27tnAqYGmOyrcs+g2xiksLchW96f1BaJ4KS
Ck61gIRRn3b4JMnXBcyxYsMZiFx6tB9hEhPcSBmtf4nSAOLHJFr6q2/JOmJhmg5y
t3ogtX4dFQmzhGfE+vi4W2YhyqmtKhORp2YtjlRstbp3mg5y2nFCpKf9n4mLV0lv
FwQpS2RjSP5jXt8TwIAq1iasENTYU60mjm9eD8dYmgetyR1/EWv+PlIawrLvqNr1
cO2z6c4vWcw6dJYJ2IFBm6lK6akAkMhRWiTfgS8p0zXWabGMi7yjAsbKiyLi2H8+
/XgY99AMM3EyjOpXNW5TgMo/zbbZXjXUnVKf6kPSkqA00oNaj5xOe9/CznQ3Mgkf
jsh6FHan9J0PwLimZYPpTtuk3s2jLgEHh44SHIOhz/0TmC8hjF2LR53rhUVet7jG
oaaR7jkqiQCHhjChC56eTco4ibHwtmiFEXLwHjlixFt7ptN+CFcm7JphSmrPmZfI
VwdIBqWHyHiYD+AsbOnxuOCjjWF2zfmiYRbLYGmCngjf8ZC51RH4DNY7TaW/5ATG
LQrLZJN47t1kA2XlVVJuRxMUIv0S54+ddNn1p4XyR5/tjcLsbv32cpx1WngJTmx2
JnyYoOPxwZQTjYHRKyFAoZM1DA9HiK2d/Ea2PycYtqGbMrah0g9KS7RwvE2CKQ70
tMCtfebkd/oQDYt7mrgLu7yve5RtW0HEJeidbey5nOtdSi8sGhRJGXINfG1U4P6N
MGiMSOfzu8ge3MbQ0d1uDgM7d5yztUAcz54V4Axr5xdKjbkgXXu6UMVttYS59xQi
zJ5uc8ne3FRBBp5dY/ACRql6NOfAkhcfeGe7EwGDrhiRcRb/REmc67Z0GDFFVgZh
SvelH15MJ+7QZc57rfLWPrApoRpXq8uUh6ptcf908AgTiV0vLuoi7rUa5A7tZJxm
XX88S0wamzSGqR1lzkmBmFwCUfN9HNx+RjA2IENlbmouPV3LGHjQzRjUElTRnIhw
MXe/4h5EwJ3TXgDQcbH+4qneVBuu5PETsnybzHPX43l0DJsADsR5OnQX0G/wB1Ez
9h8+nt7NqrcDH7qWZQsT/BbwJftJkQw3xy2hfzOvJ8G/IijDlMJV+WETENFr5r6v
DcsZUOVfiGrKzxOA4mjOjkrlQJ+BgApHBCk0vdPU1QlJDzQHYytLkKjTCVtfJ9P1
8uRd+7B6pXTgcJybPHC73vKOtarSmxJcn56CmIt3SmBa3WawITI6j8ydpV7GHVvV
/DKByM6qTiv1ha9Vo9l3o2c6erPxEcx6b+wtHWI2ZALKdVh4bZ0ZSqdZdCslks24
H0U7BGft+bl5f/Er012FQk18ILkECy+Rzy1qf0NDdzvZC+xmBtIAnKIb6cjacYQm
UFkyJ9c+eG7vjub2+V8+eqAqg0GGiHSoKfAwzGlpmD2s6+Cn16QUhuu9IPc3hyBh
iCB3jlgP4MDkplQ0uy0PJ/vfZ+sJI2sc50EJQNKdNMHyLj9HJA/ocUicrOVUROUP
cXKeTgnRJkARfzgeZiz346ENAIxK++ehUYuwufnYS8SbBqgWncVd0ciG8MmvxT+U
jUQwbxCAuWcjmffZ1zqHf1ZIElQwJ6VfGl00r/SJpQe1/2zDoiRfM2D/0y5HsPpT
0Omk59nCYUinNfZzsXYldbSbcBiXZ+W0PdA7dOIEpZh0Ft6kEvCviMxcsSDOXCp0
SW3Sid6Y3x+8xNPs26CCaQLZKWnCEv/EpSp925ofsJpIrmmgE85WHQnkopjFXTWB
G7xiLm+26nKtEZUrFMbTO1CPVGsqqj2b5ALv1UIUCtYQUZKdxsTIUdY9nXfZYt0K
qmiNLpPR/1aLTEzgg/G/fi1yOrF+3kdnpjptSK5zLmkwXANiKkoQG/2CfvB4mUrB
/M7F0bEzHi+4RQ9wXnOBgKPDY670kyyIqQYNYX2k99/ew8nm/O8E7N5ykR4fdsTh
cYps/7REM1IGT47HpkBWMul8526uH207EPI5Iu7ftA9GA6AliDtMkZH6fhyJ8faO
fKvk+0nekRHaOhA4jWFhKT2mDu+cGKW4+O3sXQa7PD0edJTE+IO4BZvpTmI5kfhF
NNQnr2pppWWrST2ajhXbx80C/dGe30qoSo7YIfYmUoTwH5ZhLCW37Q2E8qu5b6gZ
DqgirShVML+Rq/9JNbYdYStVrLzqiqnHvMFybl5dYoTfu5GuMy38YRArbi+ZkUgg
wtXYHlpuUku6mbHLdCid934JB7QRNwvNfYCkgJhsOVSICHBEjjjEM7PrtXHrYm3a
+1WBK6mkNXuh6r4ei0E0O/HGjWpH5OLxid+2GzjUtqAzZRDlTo5MUNesbkmGuXph
cxS+3FtECihFGoM5+p/GWG02lWRRHbGAMkeaXaz9mogke0TrjXf0FlIUOdx3GlRp
lsdJ3Qsc+PibJxElWVTrwJItcHMyH2K7O2e58Fg0fUvTkSvGLJ9PRPWjLHALleX1
15QfBfuyE/Y69jYF3B3762mmFNVJXZ6gk6BL6WEgD5m8KWj1Z1fMRNaJ43fzSVwu
aJnVc+LCPMwC0CyqHCKWlUqFCZh1gJjnFCKyPKK2dtH67oqZVLoh1WACPjVaO6m7
0gjLYNTFRbZ9Y4B8JFVK8IyFPj43SrS7NULEZo2uYiiy42Ec8nhrh8J7qnUsVN2W
qtRfVvmP9QKahjZGH0U6cF+/FM/K4HQrIBsJcdDIRhSq/hEX0y51kWf0oPFThHZL
L2M4/AzNAkI2PqF5hwkWJ9tMcQ+xhSVR4htrIEcgsu3AGuhFBeFKv1qe5YOkGbyE
PyhR0YqUiQlpS3eWKORk50Xb7sSoxUxe3z9C668Pwr2UmLQyC2fT9gqTSdnB/bSP
GxjIn6xSDVjh+r6YyZwqgSgSReyaOXgAn5kGI1CpNG9X187GeLPGUv4Z1DdzV5fh
BduAgA5e71DzUAMkwXvtm8IYVL1OodqC6PtrL5TzwQXCWZLdmSuyQoSFyK39VzT1
JGVjlJvWx3jM6r0bkMfib99g6PQJd8abfVsnnzklXkKA1/fHHxfzx8cIT+can41S
CZAKOV86jmOSDb56sDGf67UjdePIpRpdGLcxZ7G02O3xcGLXOF4RY1HSSizt/59Z
gld8tFeTOTA4ZN4lrv+xGApZF4eE7l0LTkMO4ISc09hEZOVhZ5bxF0mD8ZOfARJN
Q3M7R2LyzsWJ8yG0dpoLC6iFjQLRQK94Ii5LEUEDsI2Hf4+obvZIiSQ7xyxYsRVG
6bDkUp9FRtu4lAcLRNbml07f6stTm+7hdirsDEYcvCHnB2sw1T3Z/KA2Px+1BAMM
wHRZsamJBtYNsvYAQ36UqxMlf5C5Wd4gszeYoEOrWERBwOTFeY2Y8Aq+9KrlYZD6
+ODhHxnD24KXv+GJyl3LZJWAlYzfg685SbH6eZXjcVsxOKIFYgWFZTez/KKtuw0k
W9enEs7Ag54K1IJRg4iZi10/OU5754eWN4BeRJymkJv6npEs9r3jJwHOqu4ST6GC
BsK17YiG3Cug4hIMIe1AiUrKT/G+GHwaYv6V4V+k40JtWu/aw1YtW9/sg8R1Ebnl
dDbHAIWnGWBuS5XgiARi+J/Bh2srO+nC7VEtftKBn0ToedzHnX0O2s5+zrj8suU7
xkzZ4Y8LOuQhDNsl0CssJw==
`pragma protect end_protected
