// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
k8GzcZIX63NhKPadTB72GuyytMv+vwiF2euYYZUJQqnV8dZbGnfdLzPBqN6+nPvIDY+Ntv3+27sT
twAFZxi4dvud2twDAlxAWqQP+8rptszO7NLMWCK+pcYwo+d90UQGgv4dfMfzfsOg731EA66hPLGJ
QNwJS8MppO/2OsS6MTdhO4go1rhS6uc9/bWuNhV6ThQZ2ysGXKJABEJ4V0KdqePlXQLwRniLRzo1
f/XFliwxB92D6j9lDKdGl7/ckRB+VAWKxu8bBlDhlB5xYCrrgjiIgvPjE14FYDPKDt5DCLmIVicH
GX2UojFIyrfcY9xmALGHWO8vZLZc+zPScQyX2g==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 5264)
kPVr8GcJ0BNMeZXDbBtnEoy0Z+zV9cvZAOac2uYcj5csK2RLR40t/r9fuQeaKfqOjDs48vYIFeNk
lEJtEUNl4i69slU82YQL3Io0u0yrEPAWS6905H1CjMh8yHOXMj7Q7eeTWi6HqNsaxq9lBegxRXG2
uVJ0zGjIgzFpJNW0xhjLeevukjIh1T7YkpoEORjfGG6ayW0VpcP1i/u+m/xnwwaU7Tj++wl5Ja36
K03zejTbLra9fMh16WdTm0d7V3+V+MiK/Gg8BkWkJ4MWgqUUj1Lt38VrJMbitIRe9VntD2t/F4en
zMgOu5Q5Fau3ZnrQfTzXVZn/H1ezWUEk9Lg9E13S1zKYmdj9h9CKEFLv6qVaGP1czc7A+WOjjhaj
fvmJK6G5tkxVSq0AWcfs+bSubL26/NyTpZELl3kUsfkQPekw53k8JcZJ1NlXq2aBfTwbuflgOTpB
9R9TZQDvZXVZZjzSOZx0IbsYLC/IMDg9V6JHaC1rtSPXenHKhhheE43V7j2t20rXgGd8Byq9EYLo
NFunB4+gTeFpm/KJe+myn1weYiP+ncBzWs0I0WbEuD4+ty6zpQE1rQC/nvYPBfpyIROStXL/WsPr
mZzUl0Wjn4Tb02cqmE73vdkeVic2J2e02NzfD0tvVR4b6+lHX3Nffm8Dc8d0MIu2bZWBexV6bvke
hm8bZotV2T8JU0lVIw3Lr0UuGammEBowCSheWsYPcKsCWZgFLABJUWy0Bp9KoSNpEEa5BEBA/zML
0AT+owW2SAaLb+je+NatoAWAesVfrboUF+y1Cm3/RLnaZLeqxTjfHTqgJnnfAjUetFynSGbQyhV3
wVwu9v1TepAJjuuADeWLzCz3sXy1eCareK7uz6JmdoUAtn1mpADGGOKY3/nwtrsIXuHvCg5brk4W
NAE9cDBKe5d2qCqwCzqewMmDEL3YEkM/nbqrEkDmVeJyhLOicRK+b30GLLO/ytHKrPNFQk9OZsR2
jWykiX87SVbWwe366KPYIZne8oeI1gjswF+Jll75ZOL9JGdZO7EnwuQIngn4aT3OL7aAneAMIyMm
SoZnwWCrgN941TVuEDq/MDuZtZNWU0m6lX7dt8fVRXPZVrL+KLU7prYadEkJ0HQNN7mIZdjDClDZ
wcMYC2RJGAQzZ4cFoH3FwonrvAy41nJxRiA6+nVzYI3rbQAV2MhiG8cpWMpCExlc8bEtmF+d6QNk
QD2OcAZAY2X2HBxnw3czo/MC9PyxbTEJ910qCN2ApsC+mPK47soBwGh9Fh6Vsrin4132Drlz0mQy
mquA0ZBBrQFhuSBX3oJHbEM4Gaac2qvGDtqvWicVqLhAOrhr97QpJxRjiA4UW5FZS8FaQViW+A41
vCMPTAaExR0PyogMtPoHYhX02ckm1sVzGlm1DGDvgH9XTLDExR2SlXT8eRRuDb4DzziolzyWYxXb
7Qj7SQcylEjqznnQYz+w5TJhytq31JSbu35vTl0BiDv05NKcyJiBbzWN79kYeFN4nmKhfGoi42PX
SN05awITrNAqN+osKFUQ6hgnIpnr4ymLLgdlZ4IE+tY1eifKkdbVv8gW/DPyC19lDe55kUJsx5uu
KTT3au1YM+CUFvEXpnv6yztCBr8OmxXdy4zphDkZ8VM8wgJcKrDyZYJMCW2WyYvUoi0jUUAJyIIl
oFdhmyQzlAHu1QvbTD4amwxM7LQoRDOe+fpZB8zsET89rBNU/9zP1n/rVfPBr+CpOYHjY43qjre/
ESGI4qtvl8/Gv0b94qJ9raH9aUPfrq7H+wqmzLY6slCMtQZFIqPeHg0fRaKJ2C1VGZ8Nm7CTE+5k
8TbfdwSkjVTj1D7O9q7eu6vaicREZZ7teVq38bBiIG4CztwBWkccWEO8RMK4BX1RJ/ObSu2P4Woy
lB4KGl0uVhtMcM010BFKdvLmPLztz0hCd/+TNxYdShnEn/cbu98AyhRnqsUsmKkogAHk0B3xF7Gl
Efex8la5VRPJEGkkqV8fiu6hykmOBKbbn1i3EFyh6+zbMYI6jnZMWZTcP1PPhiEaZMhjToVWrWiv
Q4jkCjXXJ9BXYTgDJKMW1tyoI1ypfO5ZajYI+GtLlz3P5LAkzBTkulUbixf+JBYtQSNrQHbyoCf+
YcYkx2Sg2HXSUfEzuy/c9IyOH9c0PjHRGsrl5+AW9Ws343+a7TgWw5S+TA6cu3HaVSeuEVukgN7x
rdpTFh90ky8mIPbBQYdd3zdjZaBbGBFMSWKNMBZwUJBabEEu3n38P1b7/RrsvKDjKgeK2qHc5mN2
QvtBP+1fri28MDdpp70C4fGjxG/CPhdFf6sisBEWS0OE9YszzJce4boBQiGixYh+nxMSrZQNbRiU
KOwMpOSFIV2kmWK2nhN1daLLhiX6pB4sKRkns09XH/L5Ykvy99NruUpKZLyoKmWXzOOV3ZAi3mXq
sthp86uCkhaT6Yqs407By/zS5QMMoa9GMIvTtzWr30qSTOH3SwycittXwJdCmSH4kchPKiPRRdNg
MN3jBZKbo7wUo+568paMerIO7pxft2+o4kP2Qf46JyTiOvyKcaZW52kDlZiuRWTLVlHwHX9fRCkx
B9lMwE1+OmZKNc8iGLEO6RUyUZsvSnXf9QyQY2DY5gtZ6Z5063UGBXh704v1w/fATeeAOLcTYYxG
O0xsXgVFB3VAH678OsQzC/R3x90saWHc8NrO53+w0AOGGQZ4ftWROcyFy1OelycaX2ifJkxzpxz6
9km8wKYCERDENDc4NBT4KmXh8AG8H4iLoJdKDQ08zTrJwxitziowSsGG/4FwfuRvDrTDtl92wbvW
jj3+Rt/vhqKtALenQrC5SdGW7WMCSETOFyOdF0MlgoI5+DzE6FjDUo+ilaJEOmgmhJXvl66LEV9J
UH3l3JPjHH0o4YS4wsJduKSCEL4Qb69xveeodTuax/nWycRY8s6qXpgK55Wu+Kwu6SCzADxGYkDy
47vXzRtaARmFWLEerCOJHC3MYrjGEt0jo8tIIslvPrnI9j4P7LGpYhLXvODJ2pWXBw/8zStYdv6I
XYakmBUaFbnuYFh2DrIVQLtzyWCh+DVspIvRZwQjk0FibeLqTMYi4r4ruCEXdfhiZNGNrOjVwxS4
Xg1xl0A0XxoJ8qU75OMyxzYbFLVY6+AmiTN1uWwgMmMbngSl4g8HlB9gUNmmC+v9z5ZduuBDvI+M
lpD7c7dKQHqcV1RroZsQRHhv7phVp6Pl1r/qaAJd+dXgk0Fpiw/wEzQyFcQg9RincvbCobhY44Ry
Yl7JjKTw5eZ8BKysYUjBIQ4UdC9VD5Lj+oD/WzIXjSdnndS1cIvh+UgePZPw4TV8TyCmvmJ3X96n
qcEvLy/yt9E2tVLUzwB9oRn9WWqNjBbFP1VCCyV5inMFD/JbgtwIhknRZ23UaaZEcDv0BEF1kBty
/tWQWa0FyihJypvZNL3bYKeGfWmYZ34mu0Dj6HKYrnd/hU6m4jQp+j2b6BKPIU/8JYX0I9qOgHla
PuGUh/VC1SZ0p2l9c1wa0BLKvOQHRoGGmgVxoy4u0n6JLtUzXJhJOQ1dEIRETWi1aaGhtJuaVo9I
5ehZx2Ieu1kAxlUu4tWHkY6l4XrzgZXBFAT0Yr+f4UnZIZTk1YdDCUuOpti1T9nutfDlQpcMyyrb
BmQ+EBoSdUHaoGBCWLCffCk90PO6J5PvfTUySN5BbQoAFQz2abuTC6xlaE/ZvP+aWbf2wKYIR5EG
sIHWUSg5KU1EL8mVi95fV/3Drd2sLGpffVQX2EwQRUe/Si9dXmL6HEV3btSoMgfTGXgSfQb3yu1B
mfXw2PnjIEW/bmKb1rIauLn4kqOFvUVDfqzx3C/u39OX8aDT4/duSKZqq6ugcAMw6FMwhyTr9mxV
FX8Rqow7HfAGAfV4wGho3l+KoqbrOYScbqg5yIgtvjX7b3yT5LOrKWDjNgN7mnsg7mgPdKAsRqkX
ggJ3xNJwQ2Jh1pt1eIsyHxxUbW9572d2/1vpUOxK2xJrYwRr6z1wwnf9a1Pczh+1ICQfr1YhvAvk
6osBF8A6WYd4uC5V5NcTe7AQ0lGPcRa2gCG93z4Ks3AIsdkq2SDJkxzWHBPDA9KLM25+jIxUzy3M
9LAWT4jSSN1pZWkK+g6CNzokZqu+LqGaE7AqoWxYPkceSxi2Ci7bBhVpZmE94j/Hm09mKUAAFSxo
ux5EZ680rR6IeNTCFEtFeM93Fg4rntEkpW2moEkmirkDe8p2M9ero/6DX3Q7u+fRG6rNnktVQZId
fBVjg+Tgyjyuqpg1tgI4TgOPuoFQVjfKR/TPNeGx4tCijOKUKeHBs+Wv/VJpi2g3ylDEl/BgDdOY
rebAjibQIF1W7DQe1tNl5oFI+oVn1gZJthJ7AMcsDZ0Ygbi9qeUPoNI4memwzGNNvoxRzdgqHpQk
KKp0l90siUEfMV2vRgftnzOu3E9Tw7+s70YmZqpOoeMNrJ05pnwgWs1X6+1XRuPJSiH5NloCtkG+
odYqU7dUgEONj4rKIC4cVbwE01Y1VrTC4GeGSvapC8MRDuUM2iAuABCKBRLs4XRyzAnb7ZQRr097
S/NuEdvFiVZV56pJJFnikV0AfwRQY7xPQE9OC8wxAvccO8dc7F89z+2HLEvQaerCZZiA4MxHlgz1
V93Bmy+8t7SJHtdEYBf4tYmNu63NbNLjt0sn0sHTUMDLRwU0EU9kaJ4lScuhL8twf8Cm4U6axJHT
DRtxFZoEwYhbxdUKEnRcMTI796D/RVcL7l1Sky+pB8B5pSGahWexRm9ordIWTOIF0Sj2Fttwm8pm
lzOrMvkbX0TDp71h7Pgnu1uqXxqImAlk2820XJ0wxYwf9AbVdv42A7j5G5fzUqFY30dd/CWH6yAc
pKFE5QwGny1kee/Dgg5I5xYW5tKiBw2i+FXxK2qdGSm3D/SxRG4yyGjmoVQSNDj2qqBNuB/idE8M
MRrDWHCzKRDamcw16qgxtm23nem572F6IHiqvQyn436O/e+yTqGpd07zzxgQ87U9u4Iejset7HVP
C+aP4BzqwZNVNFuo6Lf9pSu+o13al26ifpmCzOkFgYEpj8etEJkb/3RDjpkwTzPHwXSiMMqz+RR8
g2nJTw9oDZjRVlLRUkTxo8sQMkOA2PhuIR8UsNzIqM98qboY+Wdad9rTVdm9H0v8HCRFKk7MtGs+
Nwj7vatbxgsoLAo8WNGA/EAK2inCIxETvvGR7JJAXPTFY1DGr2BJAj7OhmjFuNjL01Rn9H8gY4ST
IbK8AwWbg9ZZgZ/mKB5lZB5aIZ1Vc1UfaV9JvVEx4OLBPMzw7wi/jSn9t+JO9EUQtarv7BZAZ+t7
/ktmwoyPv4sc9rsz42Bx8drGzUM8aziP1hhJAP1CtdIiwfKNt2jDe5lgvK3g4aFTAwOmW+eV98NN
AW4pWZJwIcklnb2TDwJxBsyo8mlYvdjNZfHLvLa4RxE5vFtr73KNlXoRct4xpLZPacHFRZlJox1c
6wukG06Nvtu2s9vqXMeh3xL8cnXprPGyF1HFh0IRqy1KktmtjUUlfJzLYRF4NWc5Oy64u9SQZ1GV
wrJmSFC/NyCVBl4Tsurl1gqtacmXVpErOP+I3k7mVXszw9ZXjRzxXR4gIwpWjii3/KN67+fLJaJk
JwfrZ8nqfSduoPyKXDxtzfv4diHwTg9Wnvdy69OY4XPj2ntKrEveqmjRN+jupIU73Ck+2WVW0sWu
yyfnm/78MmT7nYv9mz79JehatM23j1Cd/hXCFveEzbP2LijCmBhFfrKB4lJJQgAaj/4onzxGfMHA
JyL+iQy4gOL6QGREMoVu+4KrVKXbh4MXMWIMHKrkuyt26iWzJrmW846fSUSr8JOGGHTN2RWxRYwE
h/aeK1T9D4f2cJ0soGLgqxe0U/v20++TUlh6ZclgWJKd8diT3HlmzuI5XRhpEFNzQmdG6zYgDocs
Puh5I3iuG4+NPkhFrPbF+wzxi+v0JSzWMCXVrv8TjM3o7uQmmglsTNRs4YXdkvfsRBpxC406a5V6
EIv/s+mXzrKfc/WZJacsoXbhLaAvhgNK1OR75TvSFNgsBPfQp31l82TC0jZEbVnzfonoJCptOWuh
m5DgSMHYhbFrzLrrdReA+8dcNvAYFNDvGNyK+g6knn56WkvrRvPuuzlSGw6Evh43z2h7P8cP139E
QKfGb+mKorP5wtTMRagU03j8SIo+ph8tdSoQ2kcYTk2I0KXrc/TO7jmm/FA+0wJF1iHZdqjJ8PAa
mSdV3cEPFR6n1U0b2V1e3gSJVaerR0giXo9ci32bPcNM6inELF9KEt4vHbm586OtALKjilT0z2kM
fX4AqbqBFqIlEtrJJcsHTkrcyw+kyCCqQ6wG5ON3xRJkk14IGOrS2a46YaFxOFHTO9X7HMONE8i9
80Ury4rkSW5JSS84Yzsrb3U8CG63A6L/PVxRaCJOx6AbqMpZmoxvfo9wd/gILNIw7/OT9y5vGvc1
1Hw5dR/M5msTj1Ee3uZMVIOX1u8ePC3qnWoyvJPlOgbDW0C+n/pv6CVkhTKfLqaq56Y4YM8MM2Vr
YFlS9CDU+kJgSKvYIaxS3yq1sYPtqjTE+BsRgQ5QDkf24rAU8mhc8URXaAr9ikVPErzlJ57XrRFl
ltlZWKp2H3eSJW5tLqmEpLGLMOlB/3KXsACCJ7cQxL87EvZmQHWvYn9jH7Ogwq2afZlyx9Ldh8j4
bwi5TfW1MgX8W9eBDVQRMU1dC4tGvKLrISyGPXlqWlqd2Y+h4tYIYcQiEv+VvH3j+1sYTBOGwyKZ
5VzmwiSVUTynF9g9LOY0AZEowNI3aSidsRB2z0KMpKj2PQLAtjkbEttWW/CTK6NUh7zNXWtmpHF/
ye994YFU0TwYzUvOXsmPrTZna4q78UGm++JOrVjU3sIHVwbfnYf0NZZ3pu5xPWZxsxZrx3RquqBD
+/R35ffWHPkLRIHKt9oDS6+b0gjzwbKJ3G4ORpCz7812hUqid2MU9aNEvLdeX8tk1dqVdWBgfuZK
Ef0picSDklJaVpC9ZsA6Uy/xctU=
`pragma protect end_protected
